
module unsaved (
	clk_clk);	

	input		clk_clk;
endmodule
