-- unsaved.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unsaved is
	port (
		clk_clk : in std_logic := '0'  -- clk.clk
	);
end entity unsaved;

architecture rtl of unsaved is
	component unsaved_buttons is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component unsaved_buttons;

	component unsaved_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(25 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(25 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component unsaved_cpu;

	component unsaved_ext_bus is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			avalon_readdata    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			avalon_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			avalon_byteenable  : out std_logic_vector(1 downto 0);                     -- byteenable
			avalon_read        : out std_logic;                                        -- read
			avalon_write       : out std_logic;                                        -- write
			avalon_writedata   : out std_logic_vector(15 downto 0);                    -- writedata
			avalon_address     : out std_logic_vector(11 downto 0);                    -- address
			address            : in  std_logic_vector(11 downto 0) := (others => 'X'); -- export
			byte_enable        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			read               : in  std_logic                     := 'X';             -- export
			write              : in  std_logic                     := 'X';             -- export
			write_data         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- export
			acknowledge        : out std_logic;                                        -- export
			read_data          : out std_logic_vector(15 downto 0)                     -- export
		);
	end component unsaved_ext_bus;

	component unsaved_flash is
		port (
			clk                 : in    std_logic                     := 'X';             -- clk
			data_cf             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			we_n                : out   std_logic;                                        -- export
			rfu                 : out   std_logic;                                        -- export
			reset_n_cf          : out   std_logic;                                        -- export
			power               : out   std_logic;                                        -- export
			iowr_n              : out   std_logic;                                        -- export
			iord_n              : out   std_logic;                                        -- export
			cs_n                : out   std_logic_vector(1 downto 0);                     -- export
			addr                : out   std_logic_vector(10 downto 0);                    -- export
			iordy               : in    std_logic                     := 'X';             -- export
			intrq               : in    std_logic                     := 'X';             -- export
			detect_n            : in    std_logic                     := 'X';             -- export
			atasel_n            : out   std_logic;                                        -- export
			av_reset_n          : in    std_logic                     := 'X';             -- reset_n
			av_ide_chipselect_n : in    std_logic                     := 'X';             -- chipselect_n
			av_ide_read_n       : in    std_logic                     := 'X';             -- read_n
			av_ide_write_n      : in    std_logic                     := 'X';             -- write_n
			av_ide_writedata    : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			av_ide_address      : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			av_ide_readdata     : out   std_logic_vector(15 downto 0);                    -- readdata
			av_ide_irq          : out   std_logic;                                        -- irq
			av_ctl_irq          : out   std_logic;                                        -- irq
			av_ctl_address      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			av_ctl_chipselect_n : in    std_logic                     := 'X';             -- chipselect_n
			av_ctl_read_n       : in    std_logic                     := 'X';             -- read_n
			av_ctl_write_n      : in    std_logic                     := 'X';             -- write_n
			av_ctl_readdata     : out   std_logic_vector(3 downto 0);                     -- readdata
			av_ctl_writedata    : in    std_logic_vector(3 downto 0)  := (others => 'X')  -- writedata
		);
	end component unsaved_flash;

	component unsaved_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component unsaved_jtag_uart_0;

	component unsaved_lcd_16207_0 is
		port (
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			clk           : in    std_logic                    := 'X';             -- clk
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic;                                       -- export
			LCD_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic                                        -- export
		);
	end component unsaved_lcd_16207_0;

	component unsaved_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component unsaved_leds;

	component unsaved_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(31 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(31 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(3 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component unsaved_sdram;

	component unsaved_sram_0 is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR     : out   std_logic_vector(19 downto 0);                    -- export
			SRAM_LB_N     : out   std_logic;                                        -- export
			SRAM_UB_N     : out   std_logic;                                        -- export
			SRAM_CE_N     : out   std_logic;                                        -- export
			SRAM_OE_N     : out   std_logic;                                        -- export
			SRAM_WE_N     : out   std_logic;                                        -- export
			address       : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			byteenable    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			read          : in    std_logic                     := 'X';             -- read
			write         : in    std_logic                     := 'X';             -- write
			writedata     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(15 downto 0);                    -- readdata
			readdatavalid : out   std_logic                                         -- readdatavalid
		);
	end component unsaved_sram_0;

	component unsaved_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component unsaved_timer_0;

	component unsaved_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component unsaved_uart_0;

	component unsaved_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			ext_bus_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			ext_bus_avalon_master_address             : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			ext_bus_avalon_master_waitrequest         : out std_logic;                                        -- waitrequest
			ext_bus_avalon_master_byteenable          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			ext_bus_avalon_master_read                : in  std_logic                     := 'X';             -- read
			ext_bus_avalon_master_readdata            : out std_logic_vector(15 downto 0);                    -- readdata
			ext_bus_avalon_master_write               : in  std_logic                     := 'X';             -- write
			ext_bus_avalon_master_writedata           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			flash_ctl_address                         : out std_logic_vector(1 downto 0);                     -- address
			flash_ctl_write                           : out std_logic;                                        -- write
			flash_ctl_read                            : out std_logic;                                        -- read
			flash_ctl_readdata                        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- readdata
			flash_ctl_writedata                       : out std_logic_vector(3 downto 0);                     -- writedata
			flash_ctl_chipselect                      : out std_logic;                                        -- chipselect
			flash_ide_address                         : out std_logic_vector(3 downto 0);                     -- address
			flash_ide_write                           : out std_logic;                                        -- write
			flash_ide_read                            : out std_logic;                                        -- read
			flash_ide_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			flash_ide_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			flash_ide_chipselect                      : out std_logic                                         -- chipselect
		);
	end component unsaved_mm_interconnect_0;

	component unsaved_mm_interconnect_1 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			cpu_reset_n_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                   : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest               : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                      : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                     : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess               : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address            : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest        : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read               : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid      : out std_logic;                                        -- readdatavalid
			buttons_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			buttons_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_address             : out std_logic_vector(8 downto 0);                     -- address
			cpu_jtag_debug_module_write               : out std_logic;                                        -- write
			cpu_jtag_debug_module_read                : out std_logic;                                        -- read
			cpu_jtag_debug_module_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_jtag_debug_module_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_jtag_debug_module_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_jtag_debug_module_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			cpu_jtag_debug_module_debugaccess         : out std_logic;                                        -- debugaccess
			jtag_uart_0_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			lcd_16207_0_control_slave_address         : out std_logic_vector(1 downto 0);                     -- address
			lcd_16207_0_control_slave_write           : out std_logic;                                        -- write
			lcd_16207_0_control_slave_read            : out std_logic;                                        -- read
			lcd_16207_0_control_slave_readdata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			lcd_16207_0_control_slave_writedata       : out std_logic_vector(7 downto 0);                     -- writedata
			lcd_16207_0_control_slave_begintransfer   : out std_logic;                                        -- begintransfer
			leds_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                             : out std_logic;                                        -- write
			leds_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                        : out std_logic;                                        -- chipselect
			sdram_s1_address                          : out std_logic_vector(21 downto 0);                    -- address
			sdram_s1_write                            : out std_logic;                                        -- write
			sdram_s1_read                             : out std_logic;                                        -- read
			sdram_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                       : out std_logic;                                        -- chipselect
			sram_0_avalon_sram_slave_address          : out std_logic_vector(19 downto 0);                    -- address
			sram_0_avalon_sram_slave_write            : out std_logic;                                        -- write
			sram_0_avalon_sram_slave_read             : out std_logic;                                        -- read
			sram_0_avalon_sram_slave_readdata         : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sram_0_avalon_sram_slave_writedata        : out std_logic_vector(15 downto 0);                    -- writedata
			sram_0_avalon_sram_slave_byteenable       : out std_logic_vector(1 downto 0);                     -- byteenable
			sram_0_avalon_sram_slave_readdatavalid    : in  std_logic                     := 'X';             -- readdatavalid
			switches_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                        : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                          : out std_logic;                                        -- write
			timer_0_s1_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                     : out std_logic;                                        -- chipselect
			uart_0_s1_address                         : out std_logic_vector(2 downto 0);                     -- address
			uart_0_s1_write                           : out std_logic;                                        -- write
			uart_0_s1_read                            : out std_logic;                                        -- read
			uart_0_s1_readdata                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			uart_0_s1_writedata                       : out std_logic_vector(15 downto 0);                    -- writedata
			uart_0_s1_begintransfer                   : out std_logic;                                        -- begintransfer
			uart_0_s1_chipselect                      : out std_logic                                         -- chipselect
		);
	end component unsaved_mm_interconnect_1;

	component unsaved_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component unsaved_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_jtag_debug_module_reset_reset                               : std_logic;                     -- cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	signal ext_bus_avalon_master_readdata                                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:ext_bus_avalon_master_readdata -> ext_bus:avalon_readdata
	signal ext_bus_avalon_master_waitrequest                               : std_logic;                     -- mm_interconnect_0:ext_bus_avalon_master_waitrequest -> ext_bus:avalon_waitrequest
	signal ext_bus_avalon_master_byteenable                                : std_logic_vector(1 downto 0);  -- ext_bus:avalon_byteenable -> mm_interconnect_0:ext_bus_avalon_master_byteenable
	signal ext_bus_avalon_master_read                                      : std_logic;                     -- ext_bus:avalon_read -> mm_interconnect_0:ext_bus_avalon_master_read
	signal ext_bus_avalon_master_address                                   : std_logic_vector(11 downto 0); -- ext_bus:avalon_address -> mm_interconnect_0:ext_bus_avalon_master_address
	signal ext_bus_avalon_master_write                                     : std_logic;                     -- ext_bus:avalon_write -> mm_interconnect_0:ext_bus_avalon_master_write
	signal ext_bus_avalon_master_writedata                                 : std_logic_vector(15 downto 0); -- ext_bus:avalon_writedata -> mm_interconnect_0:ext_bus_avalon_master_writedata
	signal mm_interconnect_0_flash_ctl_chipselect                          : std_logic;                     -- mm_interconnect_0:flash_ctl_chipselect -> mm_interconnect_0_flash_ctl_chipselect:in
	signal mm_interconnect_0_flash_ctl_readdata                            : std_logic_vector(3 downto 0);  -- flash:av_ctl_readdata -> mm_interconnect_0:flash_ctl_readdata
	signal mm_interconnect_0_flash_ctl_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:flash_ctl_address -> flash:av_ctl_address
	signal mm_interconnect_0_flash_ctl_read                                : std_logic;                     -- mm_interconnect_0:flash_ctl_read -> mm_interconnect_0_flash_ctl_read:in
	signal mm_interconnect_0_flash_ctl_write                               : std_logic;                     -- mm_interconnect_0:flash_ctl_write -> mm_interconnect_0_flash_ctl_write:in
	signal mm_interconnect_0_flash_ctl_writedata                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:flash_ctl_writedata -> flash:av_ctl_writedata
	signal mm_interconnect_0_flash_ide_chipselect                          : std_logic;                     -- mm_interconnect_0:flash_ide_chipselect -> mm_interconnect_0_flash_ide_chipselect:in
	signal mm_interconnect_0_flash_ide_readdata                            : std_logic_vector(15 downto 0); -- flash:av_ide_readdata -> mm_interconnect_0:flash_ide_readdata
	signal mm_interconnect_0_flash_ide_address                             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:flash_ide_address -> flash:av_ide_address
	signal mm_interconnect_0_flash_ide_read                                : std_logic;                     -- mm_interconnect_0:flash_ide_read -> mm_interconnect_0_flash_ide_read:in
	signal mm_interconnect_0_flash_ide_write                               : std_logic;                     -- mm_interconnect_0:flash_ide_write -> mm_interconnect_0_flash_ide_write:in
	signal mm_interconnect_0_flash_ide_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:flash_ide_writedata -> flash:av_ide_writedata
	signal cpu_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_1:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                     : std_logic;                     -- cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_1:cpu_data_master_debugaccess
	signal cpu_data_master_address                                         : std_logic_vector(25 downto 0); -- cpu:d_address -> mm_interconnect_1:cpu_data_master_address
	signal cpu_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_1:cpu_data_master_byteenable
	signal cpu_data_master_read                                            : std_logic;                     -- cpu:d_read -> mm_interconnect_1:cpu_data_master_read
	signal cpu_data_master_write                                           : std_logic;                     -- cpu:d_write -> mm_interconnect_1:cpu_data_master_write
	signal cpu_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_1:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_1:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                  : std_logic_vector(25 downto 0); -- cpu:i_address -> mm_interconnect_1:cpu_instruction_master_address
	signal cpu_instruction_master_read                                     : std_logic;                     -- cpu:i_read -> mm_interconnect_1:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_1:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_1_sram_0_avalon_sram_slave_readdata             : std_logic_vector(15 downto 0); -- sram_0:readdata -> mm_interconnect_1:sram_0_avalon_sram_slave_readdata
	signal mm_interconnect_1_sram_0_avalon_sram_slave_address              : std_logic_vector(19 downto 0); -- mm_interconnect_1:sram_0_avalon_sram_slave_address -> sram_0:address
	signal mm_interconnect_1_sram_0_avalon_sram_slave_read                 : std_logic;                     -- mm_interconnect_1:sram_0_avalon_sram_slave_read -> sram_0:read
	signal mm_interconnect_1_sram_0_avalon_sram_slave_byteenable           : std_logic_vector(1 downto 0);  -- mm_interconnect_1:sram_0_avalon_sram_slave_byteenable -> sram_0:byteenable
	signal mm_interconnect_1_sram_0_avalon_sram_slave_readdatavalid        : std_logic;                     -- sram_0:readdatavalid -> mm_interconnect_1:sram_0_avalon_sram_slave_readdatavalid
	signal mm_interconnect_1_sram_0_avalon_sram_slave_write                : std_logic;                     -- mm_interconnect_1:sram_0_avalon_sram_slave_write -> sram_0:write
	signal mm_interconnect_1_sram_0_avalon_sram_slave_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_1:sram_0_avalon_sram_slave_writedata -> sram_0:writedata
	signal mm_interconnect_1_lcd_16207_0_control_slave_readdata            : std_logic_vector(7 downto 0);  -- lcd_16207_0:readdata -> mm_interconnect_1:lcd_16207_0_control_slave_readdata
	signal mm_interconnect_1_lcd_16207_0_control_slave_address             : std_logic_vector(1 downto 0);  -- mm_interconnect_1:lcd_16207_0_control_slave_address -> lcd_16207_0:address
	signal mm_interconnect_1_lcd_16207_0_control_slave_read                : std_logic;                     -- mm_interconnect_1:lcd_16207_0_control_slave_read -> lcd_16207_0:read
	signal mm_interconnect_1_lcd_16207_0_control_slave_begintransfer       : std_logic;                     -- mm_interconnect_1:lcd_16207_0_control_slave_begintransfer -> lcd_16207_0:begintransfer
	signal mm_interconnect_1_lcd_16207_0_control_slave_write               : std_logic;                     -- mm_interconnect_1:lcd_16207_0_control_slave_write -> lcd_16207_0:write
	signal mm_interconnect_1_lcd_16207_0_control_slave_writedata           : std_logic_vector(7 downto 0);  -- mm_interconnect_1:lcd_16207_0_control_slave_writedata -> lcd_16207_0:writedata
	signal mm_interconnect_1_uart_0_s1_chipselect                          : std_logic;                     -- mm_interconnect_1:uart_0_s1_chipselect -> uart_0:chipselect
	signal mm_interconnect_1_uart_0_s1_readdata                            : std_logic_vector(15 downto 0); -- uart_0:readdata -> mm_interconnect_1:uart_0_s1_readdata
	signal mm_interconnect_1_uart_0_s1_address                             : std_logic_vector(2 downto 0);  -- mm_interconnect_1:uart_0_s1_address -> uart_0:address
	signal mm_interconnect_1_uart_0_s1_read                                : std_logic;                     -- mm_interconnect_1:uart_0_s1_read -> mm_interconnect_1_uart_0_s1_read:in
	signal mm_interconnect_1_uart_0_s1_begintransfer                       : std_logic;                     -- mm_interconnect_1:uart_0_s1_begintransfer -> uart_0:begintransfer
	signal mm_interconnect_1_uart_0_s1_write                               : std_logic;                     -- mm_interconnect_1:uart_0_s1_write -> mm_interconnect_1_uart_0_s1_write:in
	signal mm_interconnect_1_uart_0_s1_writedata                           : std_logic_vector(15 downto 0); -- mm_interconnect_1:uart_0_s1_writedata -> uart_0:writedata
	signal mm_interconnect_1_timer_0_s1_chipselect                         : std_logic;                     -- mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_1_timer_0_s1_readdata                           : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	signal mm_interconnect_1_timer_0_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_1:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_1_timer_0_s1_write                              : std_logic;                     -- mm_interconnect_1:timer_0_s1_write -> mm_interconnect_1_timer_0_s1_write:in
	signal mm_interconnect_1_timer_0_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_1_buttons_s1_readdata                           : std_logic_vector(31 downto 0); -- buttons:readdata -> mm_interconnect_1:buttons_s1_readdata
	signal mm_interconnect_1_buttons_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_1:buttons_s1_address -> buttons:address
	signal mm_interconnect_1_switches_s1_readdata                          : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_1:switches_s1_readdata
	signal mm_interconnect_1_switches_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_1:switches_s1_address -> switches:address
	signal mm_interconnect_1_leds_s1_chipselect                            : std_logic;                     -- mm_interconnect_1:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_1_leds_s1_readdata                              : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_1:leds_s1_readdata
	signal mm_interconnect_1_leds_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_1:leds_s1_address -> leds:address
	signal mm_interconnect_1_leds_s1_write                                 : std_logic;                     -- mm_interconnect_1:leds_s1_write -> mm_interconnect_1_leds_s1_write:in
	signal mm_interconnect_1_leds_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_1:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_1_sdram_s1_chipselect                           : std_logic;                     -- mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_1_sdram_s1_readdata                             : std_logic_vector(31 downto 0); -- sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	signal mm_interconnect_1_sdram_s1_waitrequest                          : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	signal mm_interconnect_1_sdram_s1_address                              : std_logic_vector(21 downto 0); -- mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_1_sdram_s1_read                                 : std_logic;                     -- mm_interconnect_1:sdram_s1_read -> mm_interconnect_1_sdram_s1_read:in
	signal mm_interconnect_1_sdram_s1_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_1:sdram_s1_byteenable -> mm_interconnect_1_sdram_s1_byteenable:in
	signal mm_interconnect_1_sdram_s1_readdatavalid                        : std_logic;                     -- sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	signal mm_interconnect_1_sdram_s1_write                                : std_logic;                     -- mm_interconnect_1:sdram_s1_write -> mm_interconnect_1_sdram_s1_write:in
	signal mm_interconnect_1_sdram_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_1_cpu_jtag_debug_module_readdata                : std_logic_vector(31 downto 0); -- cpu:jtag_debug_module_readdata -> mm_interconnect_1:cpu_jtag_debug_module_readdata
	signal mm_interconnect_1_cpu_jtag_debug_module_waitrequest             : std_logic;                     -- cpu:jtag_debug_module_waitrequest -> mm_interconnect_1:cpu_jtag_debug_module_waitrequest
	signal mm_interconnect_1_cpu_jtag_debug_module_debugaccess             : std_logic;                     -- mm_interconnect_1:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	signal mm_interconnect_1_cpu_jtag_debug_module_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_1:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	signal mm_interconnect_1_cpu_jtag_debug_module_read                    : std_logic;                     -- mm_interconnect_1:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	signal mm_interconnect_1_cpu_jtag_debug_module_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_1:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	signal mm_interconnect_1_cpu_jtag_debug_module_write                   : std_logic;                     -- mm_interconnect_1:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	signal mm_interconnect_1_cpu_jtag_debug_module_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_1:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	signal cpu_d_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:d_irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [ext_bus:reset, irq_mapper:reset, mm_interconnect_0:ext_bus_reset_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sram_0:reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_flash_ctl_chipselect_ports_inv                : std_logic;                     -- mm_interconnect_0_flash_ctl_chipselect:inv -> flash:av_ctl_chipselect_n
	signal mm_interconnect_0_flash_ctl_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_flash_ctl_read:inv -> flash:av_ctl_read_n
	signal mm_interconnect_0_flash_ctl_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_flash_ctl_write:inv -> flash:av_ctl_write_n
	signal mm_interconnect_0_flash_ide_chipselect_ports_inv                : std_logic;                     -- mm_interconnect_0_flash_ide_chipselect:inv -> flash:av_ide_chipselect_n
	signal mm_interconnect_0_flash_ide_read_ports_inv                      : std_logic;                     -- mm_interconnect_0_flash_ide_read:inv -> flash:av_ide_read_n
	signal mm_interconnect_0_flash_ide_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_flash_ide_write:inv -> flash:av_ide_write_n
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_1_uart_0_s1_read_ports_inv                      : std_logic;                     -- mm_interconnect_1_uart_0_s1_read:inv -> uart_0:read_n
	signal mm_interconnect_1_uart_0_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_1_uart_0_s1_write:inv -> uart_0:write_n
	signal mm_interconnect_1_timer_0_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_1_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_1_leds_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_1_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_1_sdram_s1_read_ports_inv                       : std_logic;                     -- mm_interconnect_1_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_1_sdram_s1_byteenable_ports_inv                 : std_logic_vector(3 downto 0);  -- mm_interconnect_1_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_1_sdram_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_1_sdram_s1_write:inv -> sdram:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [buttons:reset_n, cpu:reset_n, flash:av_reset_n, jtag_uart_0:rst_n, lcd_16207_0:reset_n, leds:reset_n, sdram:reset_n, switches:reset_n, timer_0:reset_n, uart_0:reset_n]

begin

	buttons : component unsaved_buttons
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_buttons_s1_address,     --                  s1.address
			readdata => mm_interconnect_1_buttons_s1_readdata,    --                    .readdata
			in_port  => open                                      -- external_connection.export
		);

	cpu : component unsaved_cpu
		port map (
			clk                                   => clk_clk,                                             --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,            --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_1_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_1_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_1_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_1_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_1_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_1_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_1_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_1_cpu_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                 -- custom_instruction_master.readra
		);

	ext_bus : component unsaved_ext_bus
		port map (
			clk                => clk_clk,                           --                clk.clk
			reset              => rst_controller_reset_out_reset,    --              reset.reset
			avalon_readdata    => ext_bus_avalon_master_readdata,    --      avalon_master.readdata
			avalon_waitrequest => ext_bus_avalon_master_waitrequest, --                   .waitrequest
			avalon_byteenable  => ext_bus_avalon_master_byteenable,  --                   .byteenable
			avalon_read        => ext_bus_avalon_master_read,        --                   .read
			avalon_write       => ext_bus_avalon_master_write,       --                   .write
			avalon_writedata   => ext_bus_avalon_master_writedata,   --                   .writedata
			avalon_address     => ext_bus_avalon_master_address,     --                   .address
			address            => open,                              -- external_interface.export
			byte_enable        => open,                              --                   .export
			read               => open,                              --                   .export
			write              => open,                              --                   .export
			write_data         => open,                              --                   .export
			acknowledge        => open,                              --                   .export
			read_data          => open                               --                   .export
		);

	flash : component unsaved_flash
		port map (
			clk                 => clk_clk,                                          --      clk.clk
			data_cf             => open,                                             -- external.export
			we_n                => open,                                             --         .export
			rfu                 => open,                                             --         .export
			reset_n_cf          => open,                                             --         .export
			power               => open,                                             --         .export
			iowr_n              => open,                                             --         .export
			iord_n              => open,                                             --         .export
			cs_n                => open,                                             --         .export
			addr                => open,                                             --         .export
			iordy               => open,                                             --         .export
			intrq               => open,                                             --         .export
			detect_n            => open,                                             --         .export
			atasel_n            => open,                                             --         .export
			av_reset_n          => rst_controller_reset_out_reset_ports_inv,         --    reset.reset_n
			av_ide_chipselect_n => mm_interconnect_0_flash_ide_chipselect_ports_inv, --      ide.chipselect_n
			av_ide_read_n       => mm_interconnect_0_flash_ide_read_ports_inv,       --         .read_n
			av_ide_write_n      => mm_interconnect_0_flash_ide_write_ports_inv,      --         .write_n
			av_ide_writedata    => mm_interconnect_0_flash_ide_writedata,            --         .writedata
			av_ide_address      => mm_interconnect_0_flash_ide_address,              --         .address
			av_ide_readdata     => mm_interconnect_0_flash_ide_readdata,             --         .readdata
			av_ide_irq          => open,                                             --  ide_irq.irq
			av_ctl_irq          => open,                                             --  ctl_irq.irq
			av_ctl_address      => mm_interconnect_0_flash_ctl_address,              --      ctl.address
			av_ctl_chipselect_n => mm_interconnect_0_flash_ctl_chipselect_ports_inv, --         .chipselect_n
			av_ctl_read_n       => mm_interconnect_0_flash_ctl_read_ports_inv,       --         .read_n
			av_ctl_write_n      => mm_interconnect_0_flash_ctl_write_ports_inv,      --         .write_n
			av_ctl_readdata     => mm_interconnect_0_flash_ctl_readdata,             --         .readdata
			av_ctl_writedata    => mm_interconnect_0_flash_ctl_writedata             --         .writedata
		);

	jtag_uart_0 : component unsaved_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => open                                                             --               irq.irq
		);

	lcd_16207_0 : component unsaved_lcd_16207_0
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,                  --         reset.reset_n
			clk           => clk_clk,                                                   --           clk.clk
			begintransfer => mm_interconnect_1_lcd_16207_0_control_slave_begintransfer, -- control_slave.begintransfer
			read          => mm_interconnect_1_lcd_16207_0_control_slave_read,          --              .read
			write         => mm_interconnect_1_lcd_16207_0_control_slave_write,         --              .write
			readdata      => mm_interconnect_1_lcd_16207_0_control_slave_readdata,      --              .readdata
			writedata     => mm_interconnect_1_lcd_16207_0_control_slave_writedata,     --              .writedata
			address       => mm_interconnect_1_lcd_16207_0_control_slave_address,       --              .address
			LCD_RS        => open,                                                      --      external.export
			LCD_RW        => open,                                                      --              .export
			LCD_data      => open,                                                      --              .export
			LCD_E         => open                                                       --              .export
		);

	leds : component unsaved_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_1_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_leds_s1_readdata,        --                    .readdata
			out_port   => open                                       -- external_connection.export
		);

	sdram : component unsaved_sdram
		port map (
			clk            => clk_clk,                                         --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_1_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_1_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_1_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_1_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_1_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_1_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_1_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_1_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_1_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => open,                                            --  wire.export
			zs_ba          => open,                                            --      .export
			zs_cas_n       => open,                                            --      .export
			zs_cke         => open,                                            --      .export
			zs_cs_n        => open,                                            --      .export
			zs_dq          => open,                                            --      .export
			zs_dqm         => open,                                            --      .export
			zs_ras_n       => open,                                            --      .export
			zs_we_n        => open                                             --      .export
		);

	sram_0 : component unsaved_sram_0
		port map (
			clk           => clk_clk,                                                  --                clk.clk
			reset         => rst_controller_reset_out_reset,                           --              reset.reset
			SRAM_DQ       => open,                                                     -- external_interface.export
			SRAM_ADDR     => open,                                                     --                   .export
			SRAM_LB_N     => open,                                                     --                   .export
			SRAM_UB_N     => open,                                                     --                   .export
			SRAM_CE_N     => open,                                                     --                   .export
			SRAM_OE_N     => open,                                                     --                   .export
			SRAM_WE_N     => open,                                                     --                   .export
			address       => mm_interconnect_1_sram_0_avalon_sram_slave_address,       --  avalon_sram_slave.address
			byteenable    => mm_interconnect_1_sram_0_avalon_sram_slave_byteenable,    --                   .byteenable
			read          => mm_interconnect_1_sram_0_avalon_sram_slave_read,          --                   .read
			write         => mm_interconnect_1_sram_0_avalon_sram_slave_write,         --                   .write
			writedata     => mm_interconnect_1_sram_0_avalon_sram_slave_writedata,     --                   .writedata
			readdata      => mm_interconnect_1_sram_0_avalon_sram_slave_readdata,      --                   .readdata
			readdatavalid => mm_interconnect_1_sram_0_avalon_sram_slave_readdatavalid  --                   .readdatavalid
		);

	switches : component unsaved_buttons
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_switches_s1_address,    --                  s1.address
			readdata => mm_interconnect_1_switches_s1_readdata,   --                    .readdata
			in_port  => open                                      -- external_connection.export
		);

	timer_0 : component unsaved_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_1_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_timer_0_s1_write_ports_inv, --      .write_n
			irq        => open                                          --   irq.irq
		);

	uart_0 : component unsaved_uart_0
		port map (
			clk           => clk_clk,                                     --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address       => mm_interconnect_1_uart_0_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_1_uart_0_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_1_uart_0_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_1_uart_0_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_1_uart_0_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_1_uart_0_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_1_uart_0_s1_readdata,        --                    .readdata
			rxd           => open,                                        -- external_connection.export
			txd           => open,                                        --                    .export
			irq           => open                                         --                 irq.irq
		);

	mm_interconnect_0 : component unsaved_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                --                           clk_0_clk.clk
			ext_bus_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,         -- ext_bus_reset_reset_bridge_in_reset.reset
			ext_bus_avalon_master_address             => ext_bus_avalon_master_address,          --               ext_bus_avalon_master.address
			ext_bus_avalon_master_waitrequest         => ext_bus_avalon_master_waitrequest,      --                                    .waitrequest
			ext_bus_avalon_master_byteenable          => ext_bus_avalon_master_byteenable,       --                                    .byteenable
			ext_bus_avalon_master_read                => ext_bus_avalon_master_read,             --                                    .read
			ext_bus_avalon_master_readdata            => ext_bus_avalon_master_readdata,         --                                    .readdata
			ext_bus_avalon_master_write               => ext_bus_avalon_master_write,            --                                    .write
			ext_bus_avalon_master_writedata           => ext_bus_avalon_master_writedata,        --                                    .writedata
			flash_ctl_address                         => mm_interconnect_0_flash_ctl_address,    --                           flash_ctl.address
			flash_ctl_write                           => mm_interconnect_0_flash_ctl_write,      --                                    .write
			flash_ctl_read                            => mm_interconnect_0_flash_ctl_read,       --                                    .read
			flash_ctl_readdata                        => mm_interconnect_0_flash_ctl_readdata,   --                                    .readdata
			flash_ctl_writedata                       => mm_interconnect_0_flash_ctl_writedata,  --                                    .writedata
			flash_ctl_chipselect                      => mm_interconnect_0_flash_ctl_chipselect, --                                    .chipselect
			flash_ide_address                         => mm_interconnect_0_flash_ide_address,    --                           flash_ide.address
			flash_ide_write                           => mm_interconnect_0_flash_ide_write,      --                                    .write
			flash_ide_read                            => mm_interconnect_0_flash_ide_read,       --                                    .read
			flash_ide_readdata                        => mm_interconnect_0_flash_ide_readdata,   --                                    .readdata
			flash_ide_writedata                       => mm_interconnect_0_flash_ide_writedata,  --                                    .writedata
			flash_ide_chipselect                      => mm_interconnect_0_flash_ide_chipselect  --                                    .chipselect
		);

	mm_interconnect_1 : component unsaved_mm_interconnect_1
		port map (
			clk_0_clk_clk                             => clk_clk,                                                     --                         clk_0_clk.clk
			cpu_reset_n_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                              -- cpu_reset_n_reset_bridge_in_reset.reset
			cpu_data_master_address                   => cpu_data_master_address,                                     --                   cpu_data_master.address
			cpu_data_master_waitrequest               => cpu_data_master_waitrequest,                                 --                                  .waitrequest
			cpu_data_master_byteenable                => cpu_data_master_byteenable,                                  --                                  .byteenable
			cpu_data_master_read                      => cpu_data_master_read,                                        --                                  .read
			cpu_data_master_readdata                  => cpu_data_master_readdata,                                    --                                  .readdata
			cpu_data_master_write                     => cpu_data_master_write,                                       --                                  .write
			cpu_data_master_writedata                 => cpu_data_master_writedata,                                   --                                  .writedata
			cpu_data_master_debugaccess               => cpu_data_master_debugaccess,                                 --                                  .debugaccess
			cpu_instruction_master_address            => cpu_instruction_master_address,                              --            cpu_instruction_master.address
			cpu_instruction_master_waitrequest        => cpu_instruction_master_waitrequest,                          --                                  .waitrequest
			cpu_instruction_master_read               => cpu_instruction_master_read,                                 --                                  .read
			cpu_instruction_master_readdata           => cpu_instruction_master_readdata,                             --                                  .readdata
			cpu_instruction_master_readdatavalid      => cpu_instruction_master_readdatavalid,                        --                                  .readdatavalid
			buttons_s1_address                        => mm_interconnect_1_buttons_s1_address,                        --                        buttons_s1.address
			buttons_s1_readdata                       => mm_interconnect_1_buttons_s1_readdata,                       --                                  .readdata
			cpu_jtag_debug_module_address             => mm_interconnect_1_cpu_jtag_debug_module_address,             --             cpu_jtag_debug_module.address
			cpu_jtag_debug_module_write               => mm_interconnect_1_cpu_jtag_debug_module_write,               --                                  .write
			cpu_jtag_debug_module_read                => mm_interconnect_1_cpu_jtag_debug_module_read,                --                                  .read
			cpu_jtag_debug_module_readdata            => mm_interconnect_1_cpu_jtag_debug_module_readdata,            --                                  .readdata
			cpu_jtag_debug_module_writedata           => mm_interconnect_1_cpu_jtag_debug_module_writedata,           --                                  .writedata
			cpu_jtag_debug_module_byteenable          => mm_interconnect_1_cpu_jtag_debug_module_byteenable,          --                                  .byteenable
			cpu_jtag_debug_module_waitrequest         => mm_interconnect_1_cpu_jtag_debug_module_waitrequest,         --                                  .waitrequest
			cpu_jtag_debug_module_debugaccess         => mm_interconnect_1_cpu_jtag_debug_module_debugaccess,         --                                  .debugaccess
			jtag_uart_0_avalon_jtag_slave_address     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address,     --     jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write       => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write,       --                                  .write
			jtag_uart_0_avalon_jtag_slave_read        => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read,        --                                  .read
			jtag_uart_0_avalon_jtag_slave_readdata    => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,    --                                  .readdata
			jtag_uart_0_avalon_jtag_slave_writedata   => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,   --                                  .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                  .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                  .chipselect
			lcd_16207_0_control_slave_address         => mm_interconnect_1_lcd_16207_0_control_slave_address,         --         lcd_16207_0_control_slave.address
			lcd_16207_0_control_slave_write           => mm_interconnect_1_lcd_16207_0_control_slave_write,           --                                  .write
			lcd_16207_0_control_slave_read            => mm_interconnect_1_lcd_16207_0_control_slave_read,            --                                  .read
			lcd_16207_0_control_slave_readdata        => mm_interconnect_1_lcd_16207_0_control_slave_readdata,        --                                  .readdata
			lcd_16207_0_control_slave_writedata       => mm_interconnect_1_lcd_16207_0_control_slave_writedata,       --                                  .writedata
			lcd_16207_0_control_slave_begintransfer   => mm_interconnect_1_lcd_16207_0_control_slave_begintransfer,   --                                  .begintransfer
			leds_s1_address                           => mm_interconnect_1_leds_s1_address,                           --                           leds_s1.address
			leds_s1_write                             => mm_interconnect_1_leds_s1_write,                             --                                  .write
			leds_s1_readdata                          => mm_interconnect_1_leds_s1_readdata,                          --                                  .readdata
			leds_s1_writedata                         => mm_interconnect_1_leds_s1_writedata,                         --                                  .writedata
			leds_s1_chipselect                        => mm_interconnect_1_leds_s1_chipselect,                        --                                  .chipselect
			sdram_s1_address                          => mm_interconnect_1_sdram_s1_address,                          --                          sdram_s1.address
			sdram_s1_write                            => mm_interconnect_1_sdram_s1_write,                            --                                  .write
			sdram_s1_read                             => mm_interconnect_1_sdram_s1_read,                             --                                  .read
			sdram_s1_readdata                         => mm_interconnect_1_sdram_s1_readdata,                         --                                  .readdata
			sdram_s1_writedata                        => mm_interconnect_1_sdram_s1_writedata,                        --                                  .writedata
			sdram_s1_byteenable                       => mm_interconnect_1_sdram_s1_byteenable,                       --                                  .byteenable
			sdram_s1_readdatavalid                    => mm_interconnect_1_sdram_s1_readdatavalid,                    --                                  .readdatavalid
			sdram_s1_waitrequest                      => mm_interconnect_1_sdram_s1_waitrequest,                      --                                  .waitrequest
			sdram_s1_chipselect                       => mm_interconnect_1_sdram_s1_chipselect,                       --                                  .chipselect
			sram_0_avalon_sram_slave_address          => mm_interconnect_1_sram_0_avalon_sram_slave_address,          --          sram_0_avalon_sram_slave.address
			sram_0_avalon_sram_slave_write            => mm_interconnect_1_sram_0_avalon_sram_slave_write,            --                                  .write
			sram_0_avalon_sram_slave_read             => mm_interconnect_1_sram_0_avalon_sram_slave_read,             --                                  .read
			sram_0_avalon_sram_slave_readdata         => mm_interconnect_1_sram_0_avalon_sram_slave_readdata,         --                                  .readdata
			sram_0_avalon_sram_slave_writedata        => mm_interconnect_1_sram_0_avalon_sram_slave_writedata,        --                                  .writedata
			sram_0_avalon_sram_slave_byteenable       => mm_interconnect_1_sram_0_avalon_sram_slave_byteenable,       --                                  .byteenable
			sram_0_avalon_sram_slave_readdatavalid    => mm_interconnect_1_sram_0_avalon_sram_slave_readdatavalid,    --                                  .readdatavalid
			switches_s1_address                       => mm_interconnect_1_switches_s1_address,                       --                       switches_s1.address
			switches_s1_readdata                      => mm_interconnect_1_switches_s1_readdata,                      --                                  .readdata
			timer_0_s1_address                        => mm_interconnect_1_timer_0_s1_address,                        --                        timer_0_s1.address
			timer_0_s1_write                          => mm_interconnect_1_timer_0_s1_write,                          --                                  .write
			timer_0_s1_readdata                       => mm_interconnect_1_timer_0_s1_readdata,                       --                                  .readdata
			timer_0_s1_writedata                      => mm_interconnect_1_timer_0_s1_writedata,                      --                                  .writedata
			timer_0_s1_chipselect                     => mm_interconnect_1_timer_0_s1_chipselect,                     --                                  .chipselect
			uart_0_s1_address                         => mm_interconnect_1_uart_0_s1_address,                         --                         uart_0_s1.address
			uart_0_s1_write                           => mm_interconnect_1_uart_0_s1_write,                           --                                  .write
			uart_0_s1_read                            => mm_interconnect_1_uart_0_s1_read,                            --                                  .read
			uart_0_s1_readdata                        => mm_interconnect_1_uart_0_s1_readdata,                        --                                  .readdata
			uart_0_s1_writedata                       => mm_interconnect_1_uart_0_s1_writedata,                       --                                  .writedata
			uart_0_s1_begintransfer                   => mm_interconnect_1_uart_0_s1_begintransfer,                   --                                  .begintransfer
			uart_0_s1_chipselect                      => mm_interconnect_1_uart_0_s1_chipselect                       --                                  .chipselect
		);

	irq_mapper : component unsaved_irq_mapper
		port map (
			clk        => clk_clk,                        --       clk.clk
			reset      => rst_controller_reset_out_reset, -- clk_reset.reset
			sender_irq => cpu_d_irq_irq                   --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => cpu_jtag_debug_module_reset_reset,  -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	mm_interconnect_0_flash_ctl_chipselect_ports_inv <= not mm_interconnect_0_flash_ctl_chipselect;

	mm_interconnect_0_flash_ctl_read_ports_inv <= not mm_interconnect_0_flash_ctl_read;

	mm_interconnect_0_flash_ctl_write_ports_inv <= not mm_interconnect_0_flash_ctl_write;

	mm_interconnect_0_flash_ide_chipselect_ports_inv <= not mm_interconnect_0_flash_ide_chipselect;

	mm_interconnect_0_flash_ide_read_ports_inv <= not mm_interconnect_0_flash_ide_read;

	mm_interconnect_0_flash_ide_write_ports_inv <= not mm_interconnect_0_flash_ide_write;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_1_uart_0_s1_read_ports_inv <= not mm_interconnect_1_uart_0_s1_read;

	mm_interconnect_1_uart_0_s1_write_ports_inv <= not mm_interconnect_1_uart_0_s1_write;

	mm_interconnect_1_timer_0_s1_write_ports_inv <= not mm_interconnect_1_timer_0_s1_write;

	mm_interconnect_1_leds_s1_write_ports_inv <= not mm_interconnect_1_leds_s1_write;

	mm_interconnect_1_sdram_s1_read_ports_inv <= not mm_interconnect_1_sdram_s1_read;

	mm_interconnect_1_sdram_s1_byteenable_ports_inv <= not mm_interconnect_1_sdram_s1_byteenable;

	mm_interconnect_1_sdram_s1_write_ports_inv <= not mm_interconnect_1_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of unsaved
