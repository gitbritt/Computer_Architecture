LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.STD_LOGIC_ARITH.all;
USE ieee.STD_LOGIC_UNSIGNED.all;

ENTITY mips_control IS 
	PORT( opcode				 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			funct					 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			RegDst, ALUSrc 	 : OUT STD_LOGIC;
			Jump, Jal, Jr		 : OUT STD_LOGIC;
			Beq, Bne				 : OUT STD_LOGIC;
			MemRead, MemWrite	 : OUT STD_LOGIC;
			RegWrite, MemtoReg :	OUT STD_LOGIC;
			ALUControl			 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
			);
END mips_control;

ARCHITECTURE Behavior OF mips_control IS 
	
BEGIN

	PROCESS(opcode, funct)
	BEGIN 
		CASE opcode IS 
			WHEN "000000" =>
				CASE funct IS
					WHEN "100000" =>	--ADD
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						ALUControl <= "0010";
					WHEN "100001" =>	--ADDU
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "0010";
					WHEN "100100" =>	--AND
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "0000";
					WHEN "001000" =>	--JR
						RegDst <= '0';
						ALUSrc <= '0';
						Jump <= '1';
						Jal <= '0';
						Jr <= '1';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '0';
						MemtoReg <= '0';
						AlUControl <= "0000";
					WHEN "100111" =>	--NOR
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "1100";
					WHEN "100101" =>	--OR
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "0001";
					WHEN "101010" =>	--SLT
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "0111";
					WHEN "000000" =>	--SLL
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "1000";
					WHEN "000010" =>	--SRL
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "1001";
					WHEN "000100" => --SLLV
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "1000";
					WHEN "000110" => --SRLV
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "1001";
					WHEN "100010" =>	--SUB
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "0110";
					WHEN "100011" =>	--SUBU
						RegDst <= '1';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '1';
						MemtoReg <= '0';
						AlUControl <= "0110";
					WHEN OTHERS =>
						RegDst <= '0';
						ALUSrc <= '0';
						Jump <= '0';
						Jal <= '0';
						Jr <= '0';
						Beq <= '0';
						Bne <= '0';
						MemRead <= '0';
						MemWrite <= '0';
						RegWrite <= '0';
						MemtoReg <= '0';
						AlUControl <= "0000";
					
					
				END CASE;
			WHEN "001000" =>	--ADDI
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '0';
				AlUControl <= "0010";
			WHEN "001001" =>	--ADDIU
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '0';
				AlUControl <= "0010";
			WHEN "001100" =>	--ANDI
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '0';
				AlUControl <= "0000";
			WHEN "000100" =>	--BEQ
				RegDst <= '-';
				ALUSrc <= '0';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '1';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '0';
				MemtoReg <= '0';
				AlUControl <= "0110";
			WHEN "000101" =>	--BNE
				RegDst <= '0';
				ALUSrc <= '0';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '1';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '0';
				MemtoReg <= '0';
				AlUControl <= "0110";
			WHEN "000010" =>	--J
				RegDst <= '0';
				ALUSrc <= '0';
				Jump <= '1';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '0';
				MemtoReg <= '0';
				AlUControl <= "0000";
			WHEN "000011" =>	--JAL
				RegDst <= '0';
				ALUSrc <= '0';
				Jump <= '1';
				Jal <= '1';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '0';
				AlUControl <= "0000";
			WHEN "001111" =>	--LUI
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '0';
				AlUControl <= "1101";
			WHEN "100011" =>	--LW
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '1';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '1';
				AlUControl <= "0010";
			WHEN "001101" =>	--ORI
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '0';
				AlUControl <= "0001";
			WHEN "001010" =>	--SLTI
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '1';
				MemtoReg <= '0';
				AlUControl <= "0111";
			WHEN "101011" =>	--SW
				RegDst <= '0';
				ALUSrc <= '1';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '1';
				RegWrite <= '0';
				MemtoReg <= '0';
				AlUControl <= "0010";
			WHEN OTHERS =>	--WHEN anything else
				RegDst <= '0';
				ALUSrc <= '0';
				Jump <= '0';
				Jal <= '0';
				Jr <= '0';
				Beq <= '0';
				Bne <= '0';
				MemRead <= '0';
				MemWrite <= '0';
				RegWrite <= '0';
				MemtoReg <= '0';
				AlUControl <= "0000";
				
			
			
		END CASE;
	END PROCESS;
END Behavior;